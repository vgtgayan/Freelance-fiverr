
// Bit Encodings for RV64I (look at page 126 in riscv ISA spec 2.3-draft

`define OP_JALR   7'b1100111
`define OP_THEI	  7'b0010011
`define OP_ARITH  7'b0110011
`define OP_ANDI	  7'b0010011
`define OP_LWU	  7'b0000011
`define OP_SD	  7'b0100011
`define OP_SLLI	  7'b0010011
`define OP_ADDIW  7'b0011011
`define OP_ADDW	  7'b0111011

`define FUNCT3_ARTIH_ADDI 3'b000
`define FUNCT3_ARTIH_SLTI 3'b010
`define FUNCT3_ARTIH_SLTIU 3'b011
`define FUNCT3_ARTIH_XORI 3'b100
`define FUNCT3_ARTIH_ORI 3'b110
`define FUNCT3_ARTIH_ANDI 3'b111
`define FUNCT3_ARIIH_SLLI 3'b001
`define FUNCT3_ARIIH_SRLI 3'b101
`define FUNCT3_ARITH_SRAI 3'b101
`define FUNCT3_ARTIH_ADD 3'b000
`define FUNCT3_ARTIH_SUB 3'b000
`define FUNCT3_ARTIH_SLL 3'b001
`define FUNCT3_ARTIH_SLT 3'b010
`define FUNCT3_ARTIH_SLTU 3'b011
`define FUNCT3_ARTIH_XOR 3'b100
`define FUNCT3_ARTIH_SRL 3'b101
`define FUNCT3_ARTIH_SRA 3'b101
`define FUNCT3_ARTIH_OR 3'b110
`define FUNCT3_ARTIH_AND 3'b111

`define FUNCT3_ARTIH_ADDIW 3'b000
`define FUNCT3_ARTIH_SLLIW  3'b001
`define FUNCT3_ARTIH_SRLIW  3'b101
`define FUNCT3_ARTIH_SRAIW  3'b101
`define FUNCT3_ARTIH_ADDW  3'b000
`define FUNCT3_ARTIH_SUBW  3'b000
`define FUNCT3_ARTIH_SLLW  3'b001
`define FUNCT3_ARTIH_SRLW  3'b101
`define FUNCT3_ARTIH_SAWW  3'b101

`define FUNCT7_ARTIH_ADD  7'b0000000
//`define FUNCT7 ARTIH ADD 7'b0000000
//`define FUNCT7_ARTIH_ADD 7'b0000000
`define FUNCT7_ARTIH_SUB 7'b0100000

